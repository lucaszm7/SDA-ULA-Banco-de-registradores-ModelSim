LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY multiplexador_matricial_8bits IS
	PORT (
		a, b : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END multiplexador_matricial_8bits;

ARCHITECTURE comportamente OF multiplexador_matricial_8bits IS
BEGIN

END comportamente;