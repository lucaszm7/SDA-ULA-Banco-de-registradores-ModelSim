LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY deco5to32 IS
PORT (Rd : IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		Writable : OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END deco5to32;

ARCHITECTURE comportamento OF deco5to32 IS
BEGIN

PROCESS (Rd)
		BEGIN 
			CASE Rd IS
				WHEN "00000" => Writable <= "00000000000000000000000000000001";
				WHEN "00001" => Writable <= "00000000000000000000000000000010";
				WHEN "00010" => Writable <= "00000000000000000000000000000100";
				WHEN "00011" => Writable <= "00000000000000000000000000001000";
				WHEN "00100" => Writable <= "00000000000000000000000000010000";
				WHEN "00101" => Writable <= "00000000000000000000000000100000";
				WHEN "00110" => Writable <= "00000000000000000000000001000000";
				WHEN "00111" => Writable <= "00000000000000000000000010000000";
				WHEN "01000" => Writable <= "00000000000000000000000100000000";
				WHEN "01001" => Writable <= "00000000000000000000001000000000";
				WHEN "01010" => Writable <= "00000000000000000000010000000000";
				WHEN "01011" => Writable <= "00000000000000000000100000000000";
				WHEN "01100" => Writable <= "00000000000000000001000000000000";
				WHEN "01101" => Writable <= "00000000000000000010000000000000";
				WHEN "01110" => Writable <= "00000000000000000100000000000000";
				WHEN "01111" => Writable <= "00000000000000001000000000000000";
				WHEN "10000" => Writable <= "00000000000000010000000000000000";
				WHEN "10001" => Writable <= "00000000000000100000000000000000";
				WHEN "10010" => Writable <= "00000000000001000000000000000000";
				WHEN "10011" => Writable <= "00000000000010000000000000000000";
				WHEN "10100" => Writable <= "00000000000100000000000000000000";
				WHEN "10101" => Writable <= "00000000001000000000000000000000";
				WHEN "10110" => Writable <= "00000000010000000000000000000000";
				WHEN "10111" => Writable <= "00000000100000000000000000000000";
				WHEN "11000" => Writable <= "00000001000000000000000000000000";
				WHEN "11001" => Writable <= "00000010000000000000000000000000";
				WHEN "11010" => Writable <= "00000100000000000000000000000000";
				WHEN "11011" => Writable <= "00001000000000000000000000000000";
				WHEN "11100" => Writable <= "00010000000000000000000000000000";
				WHEN "11101" => Writable <= "00100000000000000000000000000000";
				WHEN "11110" => Writable <= "01000000000000000000000000000000";
				WHEN "11111" => Writable <= "10000000000000000000000000000000";
				WHEN OTHERS  => Writable <= "00000000000000000000000000000000";
			END CASE;
		END PROCESS;
END comportamento;