LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mux9to1 IS
	PORT(
		a, b, fSoma, fSubt, colocaValorAux : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		d : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END mux9to1;

ARCHITECTURE comportamento OF mux9to1 IS

	SIGNAL A_AND_B_NOT_B : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL A_AND_B : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL A_XOR_B : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NOT_A : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL NOT_B : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
		A_AND_B_NOT_B <= (a AND b) or (NOT b);
		A_AND_B <= a AND b;
		A_XOR_B <= a XOR b;
		NOT_A <= NOT a;
		NOT_B <= NOT b;
		
		WITH FUNCT SELECT
			d <=  fSoma WHEN "000001",
					fSubt WHEN "000010",
					A_AND_B_NOT_B WHEN "000100",
					A_AND_B WHEN "001000",
					A_XOR_B WHEN "010000",
					NOT_A WHEN "100000",
					NOT_B WHEN "110000",
					colocaValorAux WHEN "100001",
					"00000000000000000000000000000000" WHEN OTHERS;
	

END comportamento;
